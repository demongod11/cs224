`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:44:36 02/23/2022 
// Design Name: 
// Module Name:    quiz2B_part2 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module quiz2B_part2(input [4:0] din, input clk, input en, input ld, input incr, output reg [4:0] q, output reg overflow);




endmodule
